// new file 
module gate_op(
  input a,b,
  output and_out
  );
  
  and(and_out,a,b);
  
 endmodule 
